module sdcard(
	input [47:0] cmd,
	input clk,send_en,rst,miso,
	output sclk,mosi,cs
	);
	
endmodule